module sin (
    input  logic        clk,
    input  logic        rst_n,
    input  logic [15:0] x,
    input  logic        start,
    output logic [15:0] result,
    output logic        done
);

logic        load_xpowertwo;
logic        init_xpowertwo;
logic        load_mult_reg;
logic        init_mult_reg;
logic        load_result;
logic        init_result;
logic        inc_counter;
logic        init_counter;
logic        sel_mult_in;
logic        co;

sin_controller controller (
    .clk(clk),
    .rst_n(rst_n),
    .start(start),
    .co(co),
    .done(done),
    .load_xpowertwo(load_xpowertwo),
    .init_xpowertwo(init_xpowertwo),
    .load_mult_reg(load_mult_reg),
    .init_mult_reg(init_mult_reg),
    .load_result(load_result),
    .init_result(init_result),
    .inc_counter(inc_counter),
    .init_counter(init_counter),
    .sel_mult_in(sel_mult_in)
);
sin_datapath datapath (
    .clk(clk),
    .rst_n(rst_n),
    .load_xpowertwo(load_xpowertwo),
    .init_xpowertwo(init_xpowertwo),
    .load_mult_reg(load_mult_reg),
    .init_mult_reg(init_mult_reg),
    .load_result(load_result),
    .init_result(init_result),
    .inc_counter(inc_counter),
    .init_counter(init_counter),
    .sel_mult_in(sel_mult_in),
    .co(co),
    .x(x),
    .result(result)
);
endmodule